typedef enum {
    {state_names}
} state_t; 

state_t present_state, next_state;
